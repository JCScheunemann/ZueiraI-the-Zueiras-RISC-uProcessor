`ifndef _my_incl_vh_
`define _my_incl_vh_
`endif

`timescale 1 ns / 1 ns

`define MEM_START_MEM_Addr 0
`define MEM_INT_MEM_Addr 2
`define MEM_INT_CH 4
`define MEM_INT_TYPE_0to3 5
`define MEM_INT_TYPE_4to7 6
`define MEM_IO_DIR_A 7
`define MEM_IO_DATA_A 8
`define MEM_IO_DIR_B 9
`define MEM_IO_DATA_B 10
`define MEM_IO_DIR_C 11
`define MEM_IO_DATA_C 12



